LIBRARY ieee;
USE ieee.std_logic_1164.ALL; 

ENTITY Conversor_binario_bcd is
	PORT (  entrada   : in  std_logic_vector(7 downto 0);
			  unidade   : out std_logic_vector(3 downto 0);
			  dezena    : out std_logic_vector(3 downto 0);
			);
END ENTITY Conversor_binario_bcd;

ARCHITECTURE arch OF Conversor_binario_bcd IS
	
BEGIN
	 			  	
	with entrada select
	unidade <=  "0000" when "00000000", --0
					"0001" when "00000001", --1
					"0010" when "00000010", --2
					"0011" when "00000011", --3
					"0100" when "00000100", --4
					"0101" when "00000101", --5
					"0110" when "00000110", --6
					"0111" when "00000111", --7
					"1000" when "00001000", --8
					"1001" when "00001001", --9
					"0000" when "00001010", --10
					"0001" when "00001011", --11
					"0010" when "00001100", --12
					"0011" when "00001101", --13
					"0100" when "00001110", --14
					"0101" when "00001111", --15
					"0110" when "00010000", --16
					"0111" when "00010001", --17
					"1000" when "00010010", --18
					"1001" when "00010011", --19
					"0000" when "00010100", --20
					"0001" when "00010101", --21
					"0010" when "00010110", --22
					"0011" when "00010111", --23
					"0100" when "00011000", --24
					"0101" when "00011001", --25
					"0110" when "00011010", --26
					"0111" when "00011011", --27
					"1000" when "00011100", --28
					"1001" when "00011101", --29
					"0000" when "00011110", --30
					"0001" when "00011111", --31
					"0010" when "00100000", --32
					"0011" when "00100001", --33
					"0100" when "00100010", --34
					"0101" when "00100011", --35
					"0110" when "00100100", --36
					"0111" when "00100101", --37
					"1000" when "00100110", --38
					"1001" when "00100111", --39
					"0000" when "00101000", --40
					"0001" when "00101001", --41
					"0010" when "00101010", --42
					"0011" when "00101011", --43
					"0100" when "00101100", --44
					"0101" when "00101101", --45
					"0110" when "00101110", --46
					"0111" when "00101111", --47
					"1000" when "00110000", --48
					"1001" when "00110001", --49
					"0000" when "00110010", --50
					"0001" when "00110011", --51
					"0010" when "00110100", --52
					"0011" when "00110101", --53
					"0100" when "00110110", --54
					"0101" when "00110111", --55
					"0110" when "00111000", --56
					"0111" when "00111001", --57
					"1000" when "00111010", --58
					"1001" when "00111011", --59
					"0000" when "00111100", --60
					"0001" when "00111101", --61
					"0010" when "00111110", --62
					"0011" when "00111111", --63
					"0100" when "01000000", --64
					"0101" when "01000001", --65
					"0110" when "01000010", --66
					"0111" when "01000011", --67
					"1000" when "01000100", --68
					"1001" when "01000101", --69
					"0000" when "01000110", --70
					"0001" when "01000111", --71
					"0010" when "01001000", --72
					"0011" when "01001001", --73
					"0100" when "01001010", --74
					"0101" when "01001011", --75
					"0110" when "01001100", --76
					"0111" when "01001101", --77
					"1000" when "01001110", --78
					"1001" when "01001111", --79
					"0000" when "01010000", --80
					"0001" when "01010001", --81
					"0010" when "01010010", --82
					"0011" when "01010011", --83
					"0100" when "01010100", --84
					"0101" when "01010101", --85
					"0110" when "01010110", --86
					"0111" when "01010111", --87
					"1000" when "01011000", --88
					"1001" when "01011001", --89
					"0000" when "01011010", --90
					"0001" when "01011011", --91
					"0010" when "01011100", --92
					"0011" when "01011101", --93
					"0100" when "01011110", --94
					"0101" when "01011111", --95
					"0110" when "01100000", --96
					"0111" when "01100001", --97
					"1000" when "01100010", --98
					"1001" when "01100011", --99
					"0000" when others;  					
					
	with entrada select
	dezena <=   "0000" when "00000000", --0
					"0000" when "00000001", --1
					"0000" when "00000010", --2
					"0000" when "00000011", --3
					"0000" when "00000100", --4
					"0000" when "00000101", --5
					"0000" when "00000110", --6
					"0000" when "00000111", --7
					"0000" when "00001000", --8
					"0000" when "00001001", --9
					"0001" when "00001010", --10
					"0001" when "00001011", --11
					"0001" when "00001100", --12
					"0001" when "00001101", --13
					"0001" when "00001110", --14
					"0001" when "00001111", --15
					"0001" when "00010000", --16
					"0001" when "00010001", --17
					"0001" when "00010010", --18
					"0001" when "00010011", --19
					"0010" when "00010100", --20
					"0010" when "00010101", --21
					"0010" when "00010110", --22
					"0010" when "00010111", --23
					"0010" when "00011000", --24
					"0010" when "00011001", --25
					"0010" when "00011010", --26
					"0010" when "00011011", --27
					"0010" when "00011100", --28
					"0010" when "00011101", --29
					"0011" when "00011110", --30
					"0011" when "00011111", --31
					"0011" when "00100000", --32
					"0011" when "00100001", --33
					"0011" when "00100010", --34
					"0011" when "00100011", --35
					"0011" when "00100100", --36
					"0011" when "00100101", --37
					"0011" when "00100110", --38
					"0011" when "00100111", --39
					"0100" when "00101000", --40
					"0100" when "00101001", --41
					"0100" when "00101010", --42
					"0100" when "00101011", --43
					"0100" when "00101100", --44
					"0100" when "00101101", --45
					"0100" when "00101110", --46
					"0100" when "00101111", --47
					"0100" when "00110000", --48
					"0100" when "00110001", --49
					"0101" when "00110010", --50
					"0101" when "00110011", --51
					"0101" when "00110100", --52
					"0101" when "00110101", --53
					"0101" when "00110110", --54
					"0101" when "00110111", --55
					"0101" when "00111000", --56
					"0101" when "00111001", --57
					"0101" when "00111010", --58
					"0101" when "00111011", --59
					"0110" when "00111100", --60
					"0110" when "00111101", --61
					"0110" when "00111110", --62
					"0110" when "00111111", --63
					"0110" when "01000000", --64
					"0110" when "01000001", --65
					"0110" when "01000010", --66
					"0110" when "01000011", --67
					"0110" when "01000100", --68
					"0110" when "01000101", --69
					"0111" when "01000110", --70
					"0111" when "01000111", --71
					"0111" when "01001000", --72
					"0111" when "01001001", --73
					"0111" when "01001010", --74
					"0111" when "01001011", --75
					"0111" when "01001100", --76
					"0111" when "01001101", --77
					"0111" when "01001110", --78
					"0111" when "01001111", --79
					"1000" when "01010000", --80
					"1000" when "01010001", --81
					"1000" when "01010010", --82
					"1000" when "01010011", --83
					"1000" when "01010100", --84
					"1000" when "01010101", --85
					"1000" when "01010110", --86
					"1000" when "01010111", --87
					"1000" when "01011000", --88
					"1000" when "01011001", --89
					"1001" when "01011010", --90
					"1001" when "01011011", --91
					"1001" when "01011100", --92
					"1001" when "01011101", --93
					"1001" when "01011110", --94
					"1001" when "01011111", --95
					"1001" when "01100000", --96
					"1001" when "01100001", --97
					"1001" when "01100010", --98
					"1001" when "01100011", --99
					"0000" when others;  
										
END ARCHITECTURE arch;
